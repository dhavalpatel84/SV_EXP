// 80bit elastic buffer design 
module tc_pcie_elastic_buffer
(
);
endmodule :tc_pcie_elastic_buffer